`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:57:52 09/08/2014 
// Design Name: 
// Module Name:    shifter 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module shifter #(parameter N=8) (
    input signed [N-1:0] IN,
    input [4:0] shamt,
    input left, input logical, 
    output [N-1:0] OUT
    );
	 
	 assign OUT = (left) ? (IN << shamt) : 
			(logical ? IN >> shamt : IN >>> shamt);

endmodule
